// area 4054*8=32000  timing 3.09
module prodtab (
    num,price,total
);

input   [3:0] num,price;
output reg  [7:0] total;

always @(*) begin
    case ({num,price})
    8'b00000000:total= 8'd0   ; //1
    8'b00000001:total= 8'd0   ; //2
    8'b00000010:total= 8'd0   ; //3
    8'b00000011:total= 8'd0   ; //4
    8'b00000100:total= 8'd0   ; //5
    8'b00000101:total= 8'd0   ; //6
    8'b00000110:total= 8'd0   ; //7
    8'b00000111:total= 8'd0   ; //8
    8'b00001000:total= 8'd0   ; //9
    8'b00001001:total= 8'd0   ; //10
    8'b00001010:total= 8'd 0   ; //11
    8'b00001011:total= 8'd 0   ; //12
    8'b00001100:total= 8'd 0   ; //13
    8'b00001101:total= 8'd 0   ; //14
    8'b00001110:total= 8'd 0   ; //15
    8'b00001111:total= 8'd 0   ; //16
    8'b00010000:total= 8'd0   ; //17
    8'b00010001:total= 8'd1   ; //18
    8'b00010010:total= 8'd2   ; //19
    8'b00010011:total= 8'd3   ; //20
    8'b00010100:total= 8'd4   ; //21
    8'b00010101:total= 8'd5   ; //22
    8'b00010110:total= 8'd6   ; //23
    8'b00010111:total= 8'd7   ; //24
    8'b00011000:total= 8'd8   ; //25
    8'b00011001:total= 8'd9   ; //26
    8'b00011010:total= 8'd 10   ; //27
    8'b00011011:total= 8'd 11   ; //28
    8'b00011100:total= 8'd 12   ; //29
    8'b00011101:total= 8'd 13   ; //30
    8'b00011110:total= 8'd 14   ; //31
    8'b00011111:total= 8'd 15   ; //32
    8'b00100000:total= 8'd0   ; //33
    8'b00100001:total= 8'd2   ; //34
    8'b00100010:total= 8'd4   ; //35
    8'b00100011:total= 8'd6   ; //36
    8'b00100100:total= 8'd8   ; //37
    8'b00100101:total= 8'd10   ; //38
    8'b00100110:total= 8'd12   ; //39
    8'b00100111:total= 8'd14   ; //40
    8'b00101000:total= 8'd16   ; //41
    8'b00101001:total= 8'd18   ; //42
    8'b00101010:total= 8'd 20   ; //43
    8'b00101011:total= 8'd 22   ; //44
    8'b00101100:total= 8'd 24   ; //45
    8'b00101101:total= 8'd 26   ; //46
    8'b00101110:total= 8'd 28   ; //47
    8'b00101111:total= 8'd 30   ; //48
    8'b00110000:total= 8'd0   ; //49
    8'b00110001:total= 8'd3   ; //50
    8'b00110010:total= 8'd6   ; //51
    8'b00110011:total= 8'd9   ; //52
    8'b00110100:total= 8'd12   ; //53
    8'b00110101:total= 8'd15   ; //54
    8'b00110110:total= 8'd18   ; //55
    8'b00110111:total= 8'd21   ; //56
    8'b00111000:total= 8'd24   ; //57
    8'b00111001:total= 8'd27   ; //58
    8'b00111010:total= 8'd 30   ; //59
    8'b00111011:total= 8'd 33   ; //60
    8'b00111100:total= 8'd 36   ; //61
    8'b00111101:total= 8'd 39   ; //62
    8'b00111110:total= 8'd 42   ; //63
    8'b00111111:total= 8'd 45   ; //64
    8'b01000000:total= 8'd0   ; //65
    8'b01000001:total= 8'd4   ; //66
    8'b01000010:total= 8'd8   ; //67
    8'b01000011:total= 8'd12   ; //68
    8'b01000100:total= 8'd16   ; //69
    8'b01000101:total= 8'd20   ; //70
    8'b01000110:total= 8'd24   ; //71
    8'b01000111:total= 8'd28   ; //72
    8'b01001000:total= 8'd32   ; //73
    8'b01001001:total= 8'd36   ; //74
    8'b01001010:total= 8'd 40   ; //75
    8'b01001011:total= 8'd 44   ; //76
    8'b01001100:total= 8'd 48   ; //77
    8'b01001101:total= 8'd 52   ; //78
    8'b01001110:total= 8'd 56   ; //79
    8'b01001111:total= 8'd 60   ; //80
    8'b01010000:total= 8'd0   ; //81
    8'b01010001:total= 8'd5   ; //82
    8'b01010010:total= 8'd10   ; //83
    8'b01010011:total= 8'd15   ; //84
    8'b01010100:total= 8'd20   ; //85
    8'b01010101:total= 8'd25   ; //86
    8'b01010110:total= 8'd30   ; //87
    8'b01010111:total= 8'd35   ; //88
    8'b01011000:total= 8'd40   ; //89
    8'b01011001:total= 8'd45   ; //90
    8'b01011010:total= 8'd 50   ; //91
    8'b01011011:total= 8'd 55   ; //92
    8'b01011100:total= 8'd 60   ; //93
    8'b01011101:total= 8'd 65   ; //94
    8'b01011110:total= 8'd 70   ; //95
    8'b01011111:total= 8'd 75   ; //96
    8'b01100000:total= 8'd0   ; //97
    8'b01100001:total= 8'd6   ; //98
    8'b01100010:total= 8'd12   ; //99
    8'b01100011:total= 8'd18   ; //100
    8'b01100100:total= 8'd24   ; //101
    8'b01100101:total= 8'd30   ; //102
    8'b01100110:total= 8'd36   ; //103
    8'b01100111:total= 8'd42   ; //104
    8'b01101000:total= 8'd48   ; //105
    8'b01101001:total= 8'd54   ; //106
    8'b01101010:total= 8'd 60   ; //107
    8'b01101011:total= 8'd 66   ; //108
    8'b01101100:total= 8'd 72   ; //109
    8'b01101101:total= 8'd 78   ; //110
    8'b01101110:total= 8'd 84   ; //111
    8'b01101111:total= 8'd 90   ; //112
    8'b01110000:total= 8'd0   ; //113
    8'b01110001:total= 8'd7   ; //114
    8'b01110010:total= 8'd14   ; //115
    8'b01110011:total= 8'd21   ; //116
    8'b01110100:total= 8'd28   ; //117
    8'b01110101:total= 8'd35   ; //118
    8'b01110110:total= 8'd42   ; //119
    8'b01110111:total= 8'd49   ; //120
    8'b01111000:total= 8'd56   ; //121
    8'b01111001:total= 8'd63   ; //122
    8'b01111010:total= 8'd 70   ; //123
    8'b01111011:total= 8'd 77   ; //124
    8'b01111100:total= 8'd 84   ; //125
    8'b01111101:total= 8'd 91   ; //126
    8'b01111110:total= 8'd 98   ; //127
    8'b01111111:total= 8'd 105   ; //128
    8'b10000000:total= 8'd0   ; //129
    8'b10000001:total= 8'd8   ; //130
    8'b10000010:total= 8'd16   ; //131
    8'b10000011:total= 8'd24   ; //132
    8'b10000100:total= 8'd32   ; //133
    8'b10000101:total= 8'd40   ; //134
    8'b10000110:total= 8'd48   ; //135
    8'b10000111:total= 8'd56   ; //136
    8'b10001000:total= 8'd64   ; //137
    8'b10001001:total= 8'd72   ; //138
    8'b10001010:total= 8'd 80   ; //139
    8'b10001011:total= 8'd 88   ; //140
    8'b10001100:total= 8'd 96   ; //141
    8'b10001101:total= 8'd 104   ; //142
    8'b10001110:total= 8'd 112   ; //143
    8'b10001111:total= 8'd 120   ; //144
    8'b10010000:total= 8'd0   ; //145
    8'b10010001:total= 8'd9   ; //146
    8'b10010010:total= 8'd18   ; //147
    8'b10010011:total= 8'd27   ; //148
    8'b10010100:total= 8'd36   ; //149
    8'b10010101:total= 8'd45   ; //150
    8'b10010110:total= 8'd54   ; //151
    8'b10010111:total= 8'd63   ; //152
    8'b10011000:total= 8'd72   ; //153
    8'b10011001:total= 8'd81   ; //154
    8'b10011010:total= 8'd90   ; //155
    8'b10011011:total= 8'd99   ; //156
    8'b10011100:total= 8'd108   ; //157
    8'b10011101:total= 8'd117   ; //158
    8'b10011110:total= 8'd126   ; //159
    8'b10011111:total= 8'd135   ; //160
    8'b10100000:total= 8'd0   ; //161
    8'b10100001:total= 8'd10   ; //162
    8'b10100010:total= 8'd20   ; //163
    8'b10100011:total= 8'd30   ; //164
    8'b10100100:total= 8'd40   ; //165
    8'b10100101:total= 8'd50   ; //166
    8'b10100110:total= 8'd60   ; //167
    8'b10100111:total= 8'd70   ; //168
    8'b10101000:total= 8'd80   ; //169
    8'b10101001:total= 8'd90   ; //170
    8'b10101010:total= 8'd 100   ; //171
    8'b10101011:total= 8'd 110   ; //172
    8'b10101100:total= 8'd 120   ; //173
    8'b10101101:total= 8'd 130   ; //174
    8'b10101110:total= 8'd 140   ; //175
    8'b10101111:total= 8'd 150   ; //176
    8'b10110000:total= 8'd0   ; //177
    8'b10110001:total= 8'd11   ; //178
    8'b10110010:total= 8'd22   ; //179
    8'b10110011:total= 8'd33   ; //180
    8'b10110100:total= 8'd44   ; //181
    8'b10110101:total= 8'd55   ; //182
    8'b10110110:total= 8'd66   ; //183
    8'b10110111:total= 8'd77   ; //184
    8'b10111000:total= 8'd88   ; //185
    8'b10111001:total= 8'd99   ; //186
    8'b10111010:total= 8'd 110   ; //187
    8'b10111011:total= 8'd 121   ; //188
    8'b10111100:total= 8'd 132   ; //189
    8'b10111101:total= 8'd 143   ; //190
    8'b10111110:total= 8'd 154   ; //191
    8'b10111111:total= 8'd 165   ; //192
    8'b11000000:total= 8'd0   ; //193
    8'b11000001:total= 8'd12   ; //194
    8'b11000010:total= 8'd24   ; //195
    8'b11000011:total= 8'd36   ; //196
    8'b11000100:total= 8'd48   ; //197
    8'b11000101:total= 8'd60   ; //198
    8'b11000110:total= 8'd72   ; //199
    8'b11000111:total= 8'd84   ; //200
    8'b11001000:total= 8'd96   ; //201
    8'b11001001:total= 8'd108   ; //202
    8'b11001010:total= 8'd 120   ; //203
    8'b11001011:total= 8'd 132   ; //204
    8'b11001100:total= 8'd 144   ; //205
    8'b11001101:total= 8'd 156   ; //206
    8'b11001110:total= 8'd 168   ; //207
    8'b11001111:total= 8'd 180   ; //208
    8'b11010000:total= 8'd0   ; //209
    8'b11010001:total= 8'd13   ; //210
    8'b11010010:total= 8'd26   ; //211
    8'b11010011:total= 8'd39   ; //212
    8'b11010100:total= 8'd52   ; //213
    8'b11010101:total= 8'd65   ; //214
    8'b11010110:total= 8'd78   ; //215
    8'b11010111:total= 8'd91   ; //216
    8'b11011000:total= 8'd104   ; //217
    8'b11011001:total= 8'd117   ; //218
    8'b11011010:total= 8'd 130   ; //219
    8'b11011011:total= 8'd 143   ; //220
    8'b11011100:total= 8'd 156   ; //221
    8'b11011101:total= 8'd 169   ; //222
    8'b11011110:total= 8'd 182   ; //223
    8'b11011111:total= 8'd 195   ; //224
    8'b11100000:total= 8'd0   ; //225
    8'b11100001:total= 8'd14   ; //226
    8'b11100010:total= 8'd28   ; //227
    8'b11100011:total= 8'd42   ; //228
    8'b11100100:total= 8'd56   ; //229
    8'b11100101:total= 8'd70   ; //230
    8'b11100110:total= 8'd84   ; //231
    8'b11100111:total= 8'd98   ; //232
    8'b11101000:total= 8'd112   ; //233
    8'b11101001:total= 8'd126   ; //234
    8'b11101010:total= 8'd 140   ; //235
    8'b11101011:total= 8'd 154   ; //236
    8'b11101100:total= 8'd 168   ; //237
    8'b11101101:total= 8'd 182   ; //238
    8'b11101110:total= 8'd 196   ; //239
    8'b11101111:total= 8'd 210   ; //240
    8'b11110000:total= 8'd0   ; //241
    8'b11110001:total= 8'd15   ; //242
    8'b11110010:total= 8'd30   ; //243
    8'b11110011:total= 8'd45   ; //244
    8'b11110100:total= 8'd60   ; //245
    8'b11110101:total= 8'd75   ; //246
    8'b11110110:total= 8'd90   ; //247
    8'b11110111:total= 8'd105   ; //248
    8'b11111000:total= 8'd120   ; //249
    8'b11111001:total= 8'd135   ; //250
    8'b11111010:total= 8'd 150   ; //251
    8'b11111011:total= 8'd 165   ; //252
    8'b11111100:total= 8'd 180   ; //253
    8'b11111101:total= 8'd 195   ; //254
    8'b11111110:total= 8'd 210   ; //255
    8'b11111111:total= 8'd 225   ; //256
    default:total=8'd0;
    endcase
end

endmodule





