//This is Bitonic Sorter.
`include "sort2.v"

// area   = 16765
// timing = 16.64
module sort_yo
(
   input  [7:0] total7, total6, total5, total4, total3, total2, total1, total0,
   output [7:0] list7, list6, list5, list4, list3, list2, list1, list0
);


//===========================================
//   level 1
//===========================================

// wire [63:0] l1out,l2out,l3out,l4out,l5out,l6out;
wire [7:0] l1 [7:0], l2 [7:0], l3 [7:0], l4 [7:0], l5 [7:0];  // 宣告五個 8x8 的 wire 陣列


b2r b2r11(.a(total7), .b(total6), .l(l1[7]), .r(l1[6]));
b2r b2r12(.a(total3), .b(total2), .l(l1[3]), .r(l1[2]));
b2l b2l11(.a(total5), .b(total4), .l(l1[5]), .r(l1[4]));
b2l b2l12(.a(total1), .b(total0), .l(l1[1]), .r(l1[0]));


//===========================================
//   level 2
//===========================================

b2r b2r21(.a(l1[7]), .b(l1[5]), .l(l2[7]), .r(l2[5]));
b2r b2r22(.a(l1[6]), .b(l1[4]), .l(l2[6]), .r(l2[4]));
b2l b2l21(.a(l1[3]), .b(l1[1]), .l(l2[3]), .r(l2[1]));
b2l b2l22(.a(l1[2]), .b(l1[0]), .l(l2[2]), .r(l2[0]));

//===========================================
//   level 3
//===========================================

b2r b2r31(.a(l2[7]), .b(l2[6]), .l(l3[7]), .r(l3[6]));
b2r b2r32(.a(l2[5]), .b(l2[4]), .l(l3[5]), .r(l3[4]));
b2l b2l31(.a(l2[3]), .b(l2[2]), .l(l3[3]), .r(l3[2]));
b2l b2l32(.a(l2[1]), .b(l2[0]), .l(l3[1]), .r(l3[0]));

//===========================================
//   level 4
//===========================================

b2r b2r41(.a(l3[7]), .b(l3[3]), .l(l4[7]), .r(l4[3]));
b2r b2r42(.a(l3[6]), .b(l3[2]), .l(l4[6]), .r(l4[2]));
b2r b2r43(.a(l3[5]), .b(l3[1]), .l(l4[5]), .r(l4[1]));
b2r b2r44(.a(l3[4]), .b(l3[0]), .l(l4[4]), .r(l4[0]));
//===========================================
//   level 5
//===========================================

b2r b2r51(.a(l4[7]), .b(l4[5]), .l(l5[7]), .r(l5[5]));
b2r b2r52(.a(l4[6]), .b(l4[4]), .l(l5[6]), .r(l5[4]));
b2r b2r53(.a(l4[3]), .b(l4[1]), .l(l5[3]), .r(l5[1]));
b2r b2r54(.a(l4[2]), .b(l4[0]), .l(l5[2]), .r(l5[0]));

//===========================================
//   level 6
//===========================================

b2r b2r61(.a(l5[7]), .b(l5[6]), .l(list0), .r(list1));
b2r b2r62(.a(l5[5]), .b(l5[4]), .l(list2), .r(list3));
b2r b2r63(.a(l5[3]), .b(l5[2]), .l(list4), .r(list5));
b2r b2r64(.a(l5[1]), .b(l5[0]), .l(list6), .r(list7));


endmodule

module b2r (
    a,b,r,l
);

input [7:0] a,b;
output [7:0] l,r;

sort2 so0( .a(a), .b(b), .big(r), .sme(l));

endmodule

module b2l (
    a,b,l,r
);

input [7:0] a,b;
output [7:0] l,r;

sort2 so0( .a(a), .b(b), .big(l), .sme(r));

endmodule